module rom (input [9:0] address, output reg [23:0] data, output [9:0] last_address);
  assign last_address = 1023;
  always @ (*) begin
    case(address)
      10'd0: data = 24'd239463;
      10'd1: data = 24'd239463;
      10'd2: data = 24'd239463;
      10'd3: data = 24'd239463;
      10'd4: data = 24'd239463;
      10'd5: data = 24'd239463;
      10'd6: data = 24'd239463;
      10'd7: data = 24'd239463;
      10'd8: data = 24'd239463;
      10'd9: data = 24'd239463;
      10'd10: data = 24'd239463;
      10'd11: data = 24'd239463;
      10'd12: data = 24'd239463;
      10'd13: data = 24'd239463;
      10'd14: data = 24'd239463;
      10'd15: data = 24'd239463;
      10'd16: data = 24'd0;
      10'd17: data = 24'd0;
      10'd18: data = 24'd0;
      10'd19: data = 24'd0;
      10'd20: data = 24'd239463;
      10'd21: data = 24'd239463;
      10'd22: data = 24'd239463;
      10'd23: data = 24'd239463;
      10'd24: data = 24'd239463;
      10'd25: data = 24'd239463;
      10'd26: data = 24'd239463;
      10'd27: data = 24'd239463;
      10'd28: data = 24'd239463;
      10'd29: data = 24'd239463;
      10'd30: data = 24'd239463;
      10'd31: data = 24'd239463;
      10'd32: data = 24'd239463;
      10'd33: data = 24'd239463;
      10'd34: data = 24'd239463;
      10'd35: data = 24'd239463;
      10'd36: data = 24'd0;
      10'd37: data = 24'd0;
      10'd38: data = 24'd0;
      10'd39: data = 24'd0;
      10'd40: data = 24'd159846;
      10'd41: data = 24'd159846;
      10'd42: data = 24'd159846;
      10'd43: data = 24'd159846;
      10'd44: data = 24'd159846;
      10'd45: data = 24'd159846;
      10'd46: data = 24'd159846;
      10'd47: data = 24'd159846;
      10'd48: data = 24'd159846;
      10'd49: data = 24'd159846;
      10'd50: data = 24'd159846;
      10'd51: data = 24'd159846;
      10'd52: data = 24'd159846;
      10'd53: data = 24'd159846;
      10'd54: data = 24'd159846;
      10'd55: data = 24'd159846;
      10'd56: data = 24'd0;
      10'd57: data = 24'd0;
      10'd58: data = 24'd0;
      10'd59: data = 24'd0;
      10'd60: data = 24'd159846;
      10'd61: data = 24'd159846;
      10'd62: data = 24'd159846;
      10'd63: data = 24'd159846;
      10'd64: data = 24'd159846;
      10'd65: data = 24'd159846;
      10'd66: data = 24'd159846;
      10'd67: data = 24'd159846;
      10'd68: data = 24'd159846;
      10'd69: data = 24'd159846;
      10'd70: data = 24'd159846;
      10'd71: data = 24'd159846;
      10'd72: data = 24'd159846;
      10'd73: data = 24'd159846;
      10'd74: data = 24'd159846;
      10'd75: data = 24'd159846;
      10'd76: data = 24'd0;
      10'd77: data = 24'd0;
      10'd78: data = 24'd0;
      10'd79: data = 24'd0;
      10'd80: data = 24'd142045;
      10'd81: data = 24'd142045;
      10'd82: data = 24'd142045;
      10'd83: data = 24'd142045;
      10'd84: data = 24'd142045;
      10'd85: data = 24'd142045;
      10'd86: data = 24'd142045;
      10'd87: data = 24'd142045;
      10'd88: data = 24'd142045;
      10'd89: data = 24'd142045;
      10'd90: data = 24'd142045;
      10'd91: data = 24'd142045;
      10'd92: data = 24'd142045;
      10'd93: data = 24'd142045;
      10'd94: data = 24'd142045;
      10'd95: data = 24'd142045;
      10'd96: data = 24'd0;
      10'd97: data = 24'd0;
      10'd98: data = 24'd0;
      10'd99: data = 24'd0;
      10'd100: data = 24'd142045;
      10'd101: data = 24'd142045;
      10'd102: data = 24'd142045;
      10'd103: data = 24'd142045;
      10'd104: data = 24'd142045;
      10'd105: data = 24'd142045;
      10'd106: data = 24'd142045;
      10'd107: data = 24'd142045;
      10'd108: data = 24'd142045;
      10'd109: data = 24'd142045;
      10'd110: data = 24'd142045;
      10'd111: data = 24'd142045;
      10'd112: data = 24'd142045;
      10'd113: data = 24'd142045;
      10'd114: data = 24'd142045;
      10'd115: data = 24'd142045;
      10'd116: data = 24'd0;
      10'd117: data = 24'd0;
      10'd118: data = 24'd0;
      10'd119: data = 24'd0;
      10'd120: data = 24'd159846;
      10'd121: data = 24'd159846;
      10'd122: data = 24'd159846;
      10'd123: data = 24'd159846;
      10'd124: data = 24'd159846;
      10'd125: data = 24'd159846;
      10'd126: data = 24'd159846;
      10'd127: data = 24'd159846;
      10'd128: data = 24'd159846;
      10'd129: data = 24'd159846;
      10'd130: data = 24'd159846;
      10'd131: data = 24'd159846;
      10'd132: data = 24'd159846;
      10'd133: data = 24'd159846;
      10'd134: data = 24'd159846;
      10'd135: data = 24'd159846;
      10'd136: data = 24'd159846;
      10'd137: data = 24'd159846;
      10'd138: data = 24'd159846;
      10'd139: data = 24'd159846;
      10'd140: data = 24'd159846;
      10'd141: data = 24'd159846;
      10'd142: data = 24'd159846;
      10'd143: data = 24'd159846;
      10'd144: data = 24'd159846;
      10'd145: data = 24'd159846;
      10'd146: data = 24'd159846;
      10'd147: data = 24'd159846;
      10'd148: data = 24'd159846;
      10'd149: data = 24'd159846;
      10'd150: data = 24'd159846;
      10'd151: data = 24'd159846;
      10'd152: data = 24'd0;
      10'd153: data = 24'd0;
      10'd154: data = 24'd0;
      10'd155: data = 24'd0;
      10'd156: data = 24'd0;
      10'd157: data = 24'd0;
      10'd158: data = 24'd0;
      10'd159: data = 24'd0;
      10'd160: data = 24'd179083;
      10'd161: data = 24'd179083;
      10'd162: data = 24'd179083;
      10'd163: data = 24'd179083;
      10'd164: data = 24'd179083;
      10'd165: data = 24'd179083;
      10'd166: data = 24'd179083;
      10'd167: data = 24'd179083;
      10'd168: data = 24'd179083;
      10'd169: data = 24'd179083;
      10'd170: data = 24'd179083;
      10'd171: data = 24'd179083;
      10'd172: data = 24'd179083;
      10'd173: data = 24'd179083;
      10'd174: data = 24'd179083;
      10'd175: data = 24'd179083;
      10'd176: data = 24'd0;
      10'd177: data = 24'd0;
      10'd178: data = 24'd0;
      10'd179: data = 24'd0;
      10'd180: data = 24'd179083;
      10'd181: data = 24'd179083;
      10'd182: data = 24'd179083;
      10'd183: data = 24'd179083;
      10'd184: data = 24'd179083;
      10'd185: data = 24'd179083;
      10'd186: data = 24'd179083;
      10'd187: data = 24'd179083;
      10'd188: data = 24'd179083;
      10'd189: data = 24'd179083;
      10'd190: data = 24'd179083;
      10'd191: data = 24'd179083;
      10'd192: data = 24'd179083;
      10'd193: data = 24'd179083;
      10'd194: data = 24'd179083;
      10'd195: data = 24'd179083;
      10'd196: data = 24'd0;
      10'd197: data = 24'd0;
      10'd198: data = 24'd0;
      10'd199: data = 24'd0;
      10'd200: data = 24'd189969;
      10'd201: data = 24'd189969;
      10'd202: data = 24'd189969;
      10'd203: data = 24'd189969;
      10'd204: data = 24'd189969;
      10'd205: data = 24'd189969;
      10'd206: data = 24'd189969;
      10'd207: data = 24'd189969;
      10'd208: data = 24'd189969;
      10'd209: data = 24'd189969;
      10'd210: data = 24'd189969;
      10'd211: data = 24'd189969;
      10'd212: data = 24'd189969;
      10'd213: data = 24'd189969;
      10'd214: data = 24'd189969;
      10'd215: data = 24'd189969;
      10'd216: data = 24'd0;
      10'd217: data = 24'd0;
      10'd218: data = 24'd0;
      10'd219: data = 24'd0;
      10'd220: data = 24'd189969;
      10'd221: data = 24'd189969;
      10'd222: data = 24'd189969;
      10'd223: data = 24'd189969;
      10'd224: data = 24'd189969;
      10'd225: data = 24'd189969;
      10'd226: data = 24'd189969;
      10'd227: data = 24'd189969;
      10'd228: data = 24'd189969;
      10'd229: data = 24'd189969;
      10'd230: data = 24'd189969;
      10'd231: data = 24'd189969;
      10'd232: data = 24'd189969;
      10'd233: data = 24'd189969;
      10'd234: data = 24'd189969;
      10'd235: data = 24'd189969;
      10'd236: data = 24'd0;
      10'd237: data = 24'd0;
      10'd238: data = 24'd0;
      10'd239: data = 24'd0;
      10'd240: data = 24'd213310;
      10'd241: data = 24'd213310;
      10'd242: data = 24'd213310;
      10'd243: data = 24'd213310;
      10'd244: data = 24'd213310;
      10'd245: data = 24'd213310;
      10'd246: data = 24'd213310;
      10'd247: data = 24'd213310;
      10'd248: data = 24'd213310;
      10'd249: data = 24'd213310;
      10'd250: data = 24'd213310;
      10'd251: data = 24'd213310;
      10'd252: data = 24'd213310;
      10'd253: data = 24'd213310;
      10'd254: data = 24'd213310;
      10'd255: data = 24'd213310;
      10'd256: data = 24'd0;
      10'd257: data = 24'd0;
      10'd258: data = 24'd0;
      10'd259: data = 24'd0;
      10'd260: data = 24'd213310;
      10'd261: data = 24'd213310;
      10'd262: data = 24'd213310;
      10'd263: data = 24'd213310;
      10'd264: data = 24'd213310;
      10'd265: data = 24'd213310;
      10'd266: data = 24'd213310;
      10'd267: data = 24'd213310;
      10'd268: data = 24'd213310;
      10'd269: data = 24'd213310;
      10'd270: data = 24'd213310;
      10'd271: data = 24'd213310;
      10'd272: data = 24'd213310;
      10'd273: data = 24'd213310;
      10'd274: data = 24'd213310;
      10'd275: data = 24'd213310;
      10'd276: data = 24'd0;
      10'd277: data = 24'd0;
      10'd278: data = 24'd0;
      10'd279: data = 24'd0;
      10'd280: data = 24'd239463;
      10'd281: data = 24'd239463;
      10'd282: data = 24'd239463;
      10'd283: data = 24'd239463;
      10'd284: data = 24'd239463;
      10'd285: data = 24'd239463;
      10'd286: data = 24'd239463;
      10'd287: data = 24'd239463;
      10'd288: data = 24'd239463;
      10'd289: data = 24'd239463;
      10'd290: data = 24'd239463;
      10'd291: data = 24'd239463;
      10'd292: data = 24'd239463;
      10'd293: data = 24'd239463;
      10'd294: data = 24'd239463;
      10'd295: data = 24'd239463;
      10'd296: data = 24'd239463;
      10'd297: data = 24'd239463;
      10'd298: data = 24'd239463;
      10'd299: data = 24'd239463;
      10'd300: data = 24'd239463;
      10'd301: data = 24'd239463;
      10'd302: data = 24'd239463;
      10'd303: data = 24'd239463;
      10'd304: data = 24'd239463;
      10'd305: data = 24'd239463;
      10'd306: data = 24'd239463;
      10'd307: data = 24'd239463;
      10'd308: data = 24'd239463;
      10'd309: data = 24'd239463;
      10'd310: data = 24'd239463;
      10'd311: data = 24'd239463;
      10'd312: data = 24'd0;
      10'd313: data = 24'd0;
      10'd314: data = 24'd0;
      10'd315: data = 24'd0;
      10'd316: data = 24'd0;
      10'd317: data = 24'd0;
      10'd318: data = 24'd0;
      10'd319: data = 24'd0;
      10'd320: data = 24'd159846;
      10'd321: data = 24'd159846;
      10'd322: data = 24'd159846;
      10'd323: data = 24'd159846;
      10'd324: data = 24'd159846;
      10'd325: data = 24'd159846;
      10'd326: data = 24'd159846;
      10'd327: data = 24'd159846;
      10'd328: data = 24'd159846;
      10'd329: data = 24'd159846;
      10'd330: data = 24'd159846;
      10'd331: data = 24'd159846;
      10'd332: data = 24'd159846;
      10'd333: data = 24'd159846;
      10'd334: data = 24'd159846;
      10'd335: data = 24'd159846;
      10'd336: data = 24'd0;
      10'd337: data = 24'd0;
      10'd338: data = 24'd0;
      10'd339: data = 24'd0;
      10'd340: data = 24'd159846;
      10'd341: data = 24'd159846;
      10'd342: data = 24'd159846;
      10'd343: data = 24'd159846;
      10'd344: data = 24'd159846;
      10'd345: data = 24'd159846;
      10'd346: data = 24'd159846;
      10'd347: data = 24'd159846;
      10'd348: data = 24'd159846;
      10'd349: data = 24'd159846;
      10'd350: data = 24'd159846;
      10'd351: data = 24'd159846;
      10'd352: data = 24'd159846;
      10'd353: data = 24'd159846;
      10'd354: data = 24'd159846;
      10'd355: data = 24'd159846;
      10'd356: data = 24'd0;
      10'd357: data = 24'd0;
      10'd358: data = 24'd0;
      10'd359: data = 24'd0;
      10'd360: data = 24'd179083;
      10'd361: data = 24'd179083;
      10'd362: data = 24'd179083;
      10'd363: data = 24'd179083;
      10'd364: data = 24'd179083;
      10'd365: data = 24'd179083;
      10'd366: data = 24'd179083;
      10'd367: data = 24'd179083;
      10'd368: data = 24'd179083;
      10'd369: data = 24'd179083;
      10'd370: data = 24'd179083;
      10'd371: data = 24'd179083;
      10'd372: data = 24'd179083;
      10'd373: data = 24'd179083;
      10'd374: data = 24'd179083;
      10'd375: data = 24'd179083;
      10'd376: data = 24'd0;
      10'd377: data = 24'd0;
      10'd378: data = 24'd0;
      10'd379: data = 24'd0;
      10'd380: data = 24'd179083;
      10'd381: data = 24'd179083;
      10'd382: data = 24'd179083;
      10'd383: data = 24'd179083;
      10'd384: data = 24'd179083;
      10'd385: data = 24'd179083;
      10'd386: data = 24'd179083;
      10'd387: data = 24'd179083;
      10'd388: data = 24'd179083;
      10'd389: data = 24'd179083;
      10'd390: data = 24'd179083;
      10'd391: data = 24'd179083;
      10'd392: data = 24'd179083;
      10'd393: data = 24'd179083;
      10'd394: data = 24'd179083;
      10'd395: data = 24'd179083;
      10'd396: data = 24'd0;
      10'd397: data = 24'd0;
      10'd398: data = 24'd0;
      10'd399: data = 24'd0;
      10'd400: data = 24'd189969;
      10'd401: data = 24'd189969;
      10'd402: data = 24'd189969;
      10'd403: data = 24'd189969;
      10'd404: data = 24'd189969;
      10'd405: data = 24'd189969;
      10'd406: data = 24'd189969;
      10'd407: data = 24'd189969;
      10'd408: data = 24'd189969;
      10'd409: data = 24'd189969;
      10'd410: data = 24'd189969;
      10'd411: data = 24'd189969;
      10'd412: data = 24'd189969;
      10'd413: data = 24'd189969;
      10'd414: data = 24'd189969;
      10'd415: data = 24'd189969;
      10'd416: data = 24'd0;
      10'd417: data = 24'd0;
      10'd418: data = 24'd0;
      10'd419: data = 24'd0;
      10'd420: data = 24'd189969;
      10'd421: data = 24'd189969;
      10'd422: data = 24'd189969;
      10'd423: data = 24'd189969;
      10'd424: data = 24'd189969;
      10'd425: data = 24'd189969;
      10'd426: data = 24'd189969;
      10'd427: data = 24'd189969;
      10'd428: data = 24'd189969;
      10'd429: data = 24'd189969;
      10'd430: data = 24'd189969;
      10'd431: data = 24'd189969;
      10'd432: data = 24'd189969;
      10'd433: data = 24'd189969;
      10'd434: data = 24'd189969;
      10'd435: data = 24'd189969;
      10'd436: data = 24'd0;
      10'd437: data = 24'd0;
      10'd438: data = 24'd0;
      10'd439: data = 24'd0;
      10'd440: data = 24'd213310;
      10'd441: data = 24'd213310;
      10'd442: data = 24'd213310;
      10'd443: data = 24'd213310;
      10'd444: data = 24'd213310;
      10'd445: data = 24'd213310;
      10'd446: data = 24'd213310;
      10'd447: data = 24'd213310;
      10'd448: data = 24'd213310;
      10'd449: data = 24'd213310;
      10'd450: data = 24'd213310;
      10'd451: data = 24'd213310;
      10'd452: data = 24'd213310;
      10'd453: data = 24'd213310;
      10'd454: data = 24'd213310;
      10'd455: data = 24'd213310;
      10'd456: data = 24'd213310;
      10'd457: data = 24'd213310;
      10'd458: data = 24'd213310;
      10'd459: data = 24'd213310;
      10'd460: data = 24'd213310;
      10'd461: data = 24'd213310;
      10'd462: data = 24'd213310;
      10'd463: data = 24'd213310;
      10'd464: data = 24'd213310;
      10'd465: data = 24'd213310;
      10'd466: data = 24'd213310;
      10'd467: data = 24'd213310;
      10'd468: data = 24'd213310;
      10'd469: data = 24'd213310;
      10'd470: data = 24'd213310;
      10'd471: data = 24'd213310;
      10'd472: data = 24'd0;
      10'd473: data = 24'd0;
      10'd474: data = 24'd0;
      10'd475: data = 24'd0;
      10'd476: data = 24'd0;
      10'd477: data = 24'd0;
      10'd478: data = 24'd0;
      10'd479: data = 24'd0;
      10'd480: data = 24'd159846;
      10'd481: data = 24'd159846;
      10'd482: data = 24'd159846;
      10'd483: data = 24'd159846;
      10'd484: data = 24'd159846;
      10'd485: data = 24'd159846;
      10'd486: data = 24'd159846;
      10'd487: data = 24'd159846;
      10'd488: data = 24'd159846;
      10'd489: data = 24'd159846;
      10'd490: data = 24'd159846;
      10'd491: data = 24'd159846;
      10'd492: data = 24'd159846;
      10'd493: data = 24'd159846;
      10'd494: data = 24'd159846;
      10'd495: data = 24'd159846;
      10'd496: data = 24'd0;
      10'd497: data = 24'd0;
      10'd498: data = 24'd0;
      10'd499: data = 24'd0;
      10'd500: data = 24'd159846;
      10'd501: data = 24'd159846;
      10'd502: data = 24'd159846;
      10'd503: data = 24'd159846;
      10'd504: data = 24'd159846;
      10'd505: data = 24'd159846;
      10'd506: data = 24'd159846;
      10'd507: data = 24'd159846;
      10'd508: data = 24'd159846;
      10'd509: data = 24'd159846;
      10'd510: data = 24'd159846;
      10'd511: data = 24'd159846;
      10'd512: data = 24'd159846;
      10'd513: data = 24'd159846;
      10'd514: data = 24'd159846;
      10'd515: data = 24'd159846;
      10'd516: data = 24'd0;
      10'd517: data = 24'd0;
      10'd518: data = 24'd0;
      10'd519: data = 24'd0;
      10'd520: data = 24'd179083;
      10'd521: data = 24'd179083;
      10'd522: data = 24'd179083;
      10'd523: data = 24'd179083;
      10'd524: data = 24'd179083;
      10'd525: data = 24'd179083;
      10'd526: data = 24'd179083;
      10'd527: data = 24'd179083;
      10'd528: data = 24'd179083;
      10'd529: data = 24'd179083;
      10'd530: data = 24'd179083;
      10'd531: data = 24'd179083;
      10'd532: data = 24'd179083;
      10'd533: data = 24'd179083;
      10'd534: data = 24'd179083;
      10'd535: data = 24'd179083;
      10'd536: data = 24'd0;
      10'd537: data = 24'd0;
      10'd538: data = 24'd0;
      10'd539: data = 24'd0;
      10'd540: data = 24'd179083;
      10'd541: data = 24'd179083;
      10'd542: data = 24'd179083;
      10'd543: data = 24'd179083;
      10'd544: data = 24'd179083;
      10'd545: data = 24'd179083;
      10'd546: data = 24'd179083;
      10'd547: data = 24'd179083;
      10'd548: data = 24'd179083;
      10'd549: data = 24'd179083;
      10'd550: data = 24'd179083;
      10'd551: data = 24'd179083;
      10'd552: data = 24'd179083;
      10'd553: data = 24'd179083;
      10'd554: data = 24'd179083;
      10'd555: data = 24'd179083;
      10'd556: data = 24'd0;
      10'd557: data = 24'd0;
      10'd558: data = 24'd0;
      10'd559: data = 24'd0;
      10'd560: data = 24'd189969;
      10'd561: data = 24'd189969;
      10'd562: data = 24'd189969;
      10'd563: data = 24'd189969;
      10'd564: data = 24'd189969;
      10'd565: data = 24'd189969;
      10'd566: data = 24'd189969;
      10'd567: data = 24'd189969;
      10'd568: data = 24'd189969;
      10'd569: data = 24'd189969;
      10'd570: data = 24'd189969;
      10'd571: data = 24'd189969;
      10'd572: data = 24'd189969;
      10'd573: data = 24'd189969;
      10'd574: data = 24'd189969;
      10'd575: data = 24'd189969;
      10'd576: data = 24'd0;
      10'd577: data = 24'd0;
      10'd578: data = 24'd0;
      10'd579: data = 24'd0;
      10'd580: data = 24'd189969;
      10'd581: data = 24'd189969;
      10'd582: data = 24'd189969;
      10'd583: data = 24'd189969;
      10'd584: data = 24'd189969;
      10'd585: data = 24'd189969;
      10'd586: data = 24'd189969;
      10'd587: data = 24'd189969;
      10'd588: data = 24'd189969;
      10'd589: data = 24'd189969;
      10'd590: data = 24'd189969;
      10'd591: data = 24'd189969;
      10'd592: data = 24'd189969;
      10'd593: data = 24'd189969;
      10'd594: data = 24'd189969;
      10'd595: data = 24'd189969;
      10'd596: data = 24'd0;
      10'd597: data = 24'd0;
      10'd598: data = 24'd0;
      10'd599: data = 24'd0;
      10'd600: data = 24'd213310;
      10'd601: data = 24'd213310;
      10'd602: data = 24'd213310;
      10'd603: data = 24'd213310;
      10'd604: data = 24'd213310;
      10'd605: data = 24'd213310;
      10'd606: data = 24'd213310;
      10'd607: data = 24'd213310;
      10'd608: data = 24'd213310;
      10'd609: data = 24'd213310;
      10'd610: data = 24'd213310;
      10'd611: data = 24'd213310;
      10'd612: data = 24'd213310;
      10'd613: data = 24'd213310;
      10'd614: data = 24'd213310;
      10'd615: data = 24'd213310;
      10'd616: data = 24'd213310;
      10'd617: data = 24'd213310;
      10'd618: data = 24'd213310;
      10'd619: data = 24'd213310;
      10'd620: data = 24'd213310;
      10'd621: data = 24'd213310;
      10'd622: data = 24'd213310;
      10'd623: data = 24'd213310;
      10'd624: data = 24'd213310;
      10'd625: data = 24'd213310;
      10'd626: data = 24'd213310;
      10'd627: data = 24'd213310;
      10'd628: data = 24'd213310;
      10'd629: data = 24'd213310;
      10'd630: data = 24'd213310;
      10'd631: data = 24'd213310;
      10'd632: data = 24'd0;
      10'd633: data = 24'd0;
      10'd634: data = 24'd0;
      10'd635: data = 24'd0;
      10'd636: data = 24'd0;
      10'd637: data = 24'd0;
      10'd638: data = 24'd0;
      10'd639: data = 24'd0;
      10'd640: data = 24'd239463;
      10'd641: data = 24'd239463;
      10'd642: data = 24'd239463;
      10'd643: data = 24'd239463;
      10'd644: data = 24'd239463;
      10'd645: data = 24'd239463;
      10'd646: data = 24'd239463;
      10'd647: data = 24'd239463;
      10'd648: data = 24'd239463;
      10'd649: data = 24'd239463;
      10'd650: data = 24'd239463;
      10'd651: data = 24'd239463;
      10'd652: data = 24'd239463;
      10'd653: data = 24'd239463;
      10'd654: data = 24'd239463;
      10'd655: data = 24'd239463;
      10'd656: data = 24'd0;
      10'd657: data = 24'd0;
      10'd658: data = 24'd0;
      10'd659: data = 24'd0;
      10'd660: data = 24'd239463;
      10'd661: data = 24'd239463;
      10'd662: data = 24'd239463;
      10'd663: data = 24'd239463;
      10'd664: data = 24'd239463;
      10'd665: data = 24'd239463;
      10'd666: data = 24'd239463;
      10'd667: data = 24'd239463;
      10'd668: data = 24'd239463;
      10'd669: data = 24'd239463;
      10'd670: data = 24'd239463;
      10'd671: data = 24'd239463;
      10'd672: data = 24'd239463;
      10'd673: data = 24'd239463;
      10'd674: data = 24'd239463;
      10'd675: data = 24'd239463;
      10'd676: data = 24'd0;
      10'd677: data = 24'd0;
      10'd678: data = 24'd0;
      10'd679: data = 24'd0;
      10'd680: data = 24'd159846;
      10'd681: data = 24'd159846;
      10'd682: data = 24'd159846;
      10'd683: data = 24'd159846;
      10'd684: data = 24'd159846;
      10'd685: data = 24'd159846;
      10'd686: data = 24'd159846;
      10'd687: data = 24'd159846;
      10'd688: data = 24'd159846;
      10'd689: data = 24'd159846;
      10'd690: data = 24'd159846;
      10'd691: data = 24'd159846;
      10'd692: data = 24'd159846;
      10'd693: data = 24'd159846;
      10'd694: data = 24'd159846;
      10'd695: data = 24'd159846;
      10'd696: data = 24'd0;
      10'd697: data = 24'd0;
      10'd698: data = 24'd0;
      10'd699: data = 24'd0;
      10'd700: data = 24'd159846;
      10'd701: data = 24'd159846;
      10'd702: data = 24'd159846;
      10'd703: data = 24'd159846;
      10'd704: data = 24'd159846;
      10'd705: data = 24'd159846;
      10'd706: data = 24'd159846;
      10'd707: data = 24'd159846;
      10'd708: data = 24'd159846;
      10'd709: data = 24'd159846;
      10'd710: data = 24'd159846;
      10'd711: data = 24'd159846;
      10'd712: data = 24'd159846;
      10'd713: data = 24'd159846;
      10'd714: data = 24'd159846;
      10'd715: data = 24'd159846;
      10'd716: data = 24'd0;
      10'd717: data = 24'd0;
      10'd718: data = 24'd0;
      10'd719: data = 24'd0;
      10'd720: data = 24'd142045;
      10'd721: data = 24'd142045;
      10'd722: data = 24'd142045;
      10'd723: data = 24'd142045;
      10'd724: data = 24'd142045;
      10'd725: data = 24'd142045;
      10'd726: data = 24'd142045;
      10'd727: data = 24'd142045;
      10'd728: data = 24'd142045;
      10'd729: data = 24'd142045;
      10'd730: data = 24'd142045;
      10'd731: data = 24'd142045;
      10'd732: data = 24'd142045;
      10'd733: data = 24'd142045;
      10'd734: data = 24'd142045;
      10'd735: data = 24'd142045;
      10'd736: data = 24'd0;
      10'd737: data = 24'd0;
      10'd738: data = 24'd0;
      10'd739: data = 24'd0;
      10'd740: data = 24'd142045;
      10'd741: data = 24'd142045;
      10'd742: data = 24'd142045;
      10'd743: data = 24'd142045;
      10'd744: data = 24'd142045;
      10'd745: data = 24'd142045;
      10'd746: data = 24'd142045;
      10'd747: data = 24'd142045;
      10'd748: data = 24'd142045;
      10'd749: data = 24'd142045;
      10'd750: data = 24'd142045;
      10'd751: data = 24'd142045;
      10'd752: data = 24'd142045;
      10'd753: data = 24'd142045;
      10'd754: data = 24'd142045;
      10'd755: data = 24'd142045;
      10'd756: data = 24'd0;
      10'd757: data = 24'd0;
      10'd758: data = 24'd0;
      10'd759: data = 24'd0;
      10'd760: data = 24'd159846;
      10'd761: data = 24'd159846;
      10'd762: data = 24'd159846;
      10'd763: data = 24'd159846;
      10'd764: data = 24'd159846;
      10'd765: data = 24'd159846;
      10'd766: data = 24'd159846;
      10'd767: data = 24'd159846;
      10'd768: data = 24'd159846;
      10'd769: data = 24'd159846;
      10'd770: data = 24'd159846;
      10'd771: data = 24'd159846;
      10'd772: data = 24'd159846;
      10'd773: data = 24'd159846;
      10'd774: data = 24'd159846;
      10'd775: data = 24'd159846;
      10'd776: data = 24'd159846;
      10'd777: data = 24'd159846;
      10'd778: data = 24'd159846;
      10'd779: data = 24'd159846;
      10'd780: data = 24'd159846;
      10'd781: data = 24'd159846;
      10'd782: data = 24'd159846;
      10'd783: data = 24'd159846;
      10'd784: data = 24'd159846;
      10'd785: data = 24'd159846;
      10'd786: data = 24'd159846;
      10'd787: data = 24'd159846;
      10'd788: data = 24'd159846;
      10'd789: data = 24'd159846;
      10'd790: data = 24'd159846;
      10'd791: data = 24'd159846;
      10'd792: data = 24'd0;
      10'd793: data = 24'd0;
      10'd794: data = 24'd0;
      10'd795: data = 24'd0;
      10'd796: data = 24'd0;
      10'd797: data = 24'd0;
      10'd798: data = 24'd0;
      10'd799: data = 24'd0;
      10'd800: data = 24'd179083;
      10'd801: data = 24'd179083;
      10'd802: data = 24'd179083;
      10'd803: data = 24'd179083;
      10'd804: data = 24'd179083;
      10'd805: data = 24'd179083;
      10'd806: data = 24'd179083;
      10'd807: data = 24'd179083;
      10'd808: data = 24'd179083;
      10'd809: data = 24'd179083;
      10'd810: data = 24'd179083;
      10'd811: data = 24'd179083;
      10'd812: data = 24'd179083;
      10'd813: data = 24'd179083;
      10'd814: data = 24'd179083;
      10'd815: data = 24'd179083;
      10'd816: data = 24'd0;
      10'd817: data = 24'd0;
      10'd818: data = 24'd0;
      10'd819: data = 24'd0;
      10'd820: data = 24'd179083;
      10'd821: data = 24'd179083;
      10'd822: data = 24'd179083;
      10'd823: data = 24'd179083;
      10'd824: data = 24'd179083;
      10'd825: data = 24'd179083;
      10'd826: data = 24'd179083;
      10'd827: data = 24'd179083;
      10'd828: data = 24'd179083;
      10'd829: data = 24'd179083;
      10'd830: data = 24'd179083;
      10'd831: data = 24'd179083;
      10'd832: data = 24'd179083;
      10'd833: data = 24'd179083;
      10'd834: data = 24'd179083;
      10'd835: data = 24'd179083;
      10'd836: data = 24'd0;
      10'd837: data = 24'd0;
      10'd838: data = 24'd0;
      10'd839: data = 24'd0;
      10'd840: data = 24'd189969;
      10'd841: data = 24'd189969;
      10'd842: data = 24'd189969;
      10'd843: data = 24'd189969;
      10'd844: data = 24'd189969;
      10'd845: data = 24'd189969;
      10'd846: data = 24'd189969;
      10'd847: data = 24'd189969;
      10'd848: data = 24'd189969;
      10'd849: data = 24'd189969;
      10'd850: data = 24'd189969;
      10'd851: data = 24'd189969;
      10'd852: data = 24'd189969;
      10'd853: data = 24'd189969;
      10'd854: data = 24'd189969;
      10'd855: data = 24'd189969;
      10'd856: data = 24'd0;
      10'd857: data = 24'd0;
      10'd858: data = 24'd0;
      10'd859: data = 24'd0;
      10'd860: data = 24'd189969;
      10'd861: data = 24'd189969;
      10'd862: data = 24'd189969;
      10'd863: data = 24'd189969;
      10'd864: data = 24'd189969;
      10'd865: data = 24'd189969;
      10'd866: data = 24'd189969;
      10'd867: data = 24'd189969;
      10'd868: data = 24'd189969;
      10'd869: data = 24'd189969;
      10'd870: data = 24'd189969;
      10'd871: data = 24'd189969;
      10'd872: data = 24'd189969;
      10'd873: data = 24'd189969;
      10'd874: data = 24'd189969;
      10'd875: data = 24'd189969;
      10'd876: data = 24'd0;
      10'd877: data = 24'd0;
      10'd878: data = 24'd0;
      10'd879: data = 24'd0;
      10'd880: data = 24'd213310;
      10'd881: data = 24'd213310;
      10'd882: data = 24'd213310;
      10'd883: data = 24'd213310;
      10'd884: data = 24'd213310;
      10'd885: data = 24'd213310;
      10'd886: data = 24'd213310;
      10'd887: data = 24'd213310;
      10'd888: data = 24'd213310;
      10'd889: data = 24'd213310;
      10'd890: data = 24'd213310;
      10'd891: data = 24'd213310;
      10'd892: data = 24'd213310;
      10'd893: data = 24'd213310;
      10'd894: data = 24'd213310;
      10'd895: data = 24'd213310;
      10'd896: data = 24'd0;
      10'd897: data = 24'd0;
      10'd898: data = 24'd0;
      10'd899: data = 24'd0;
      10'd900: data = 24'd213310;
      10'd901: data = 24'd213310;
      10'd902: data = 24'd213310;
      10'd903: data = 24'd213310;
      10'd904: data = 24'd213310;
      10'd905: data = 24'd213310;
      10'd906: data = 24'd213310;
      10'd907: data = 24'd213310;
      10'd908: data = 24'd213310;
      10'd909: data = 24'd213310;
      10'd910: data = 24'd213310;
      10'd911: data = 24'd213310;
      10'd912: data = 24'd213310;
      10'd913: data = 24'd213310;
      10'd914: data = 24'd213310;
      10'd915: data = 24'd213310;
      10'd916: data = 24'd0;
      10'd917: data = 24'd0;
      10'd918: data = 24'd0;
      10'd919: data = 24'd0;
      10'd920: data = 24'd239463;
      10'd921: data = 24'd239463;
      10'd922: data = 24'd239463;
      10'd923: data = 24'd239463;
      10'd924: data = 24'd239463;
      10'd925: data = 24'd239463;
      10'd926: data = 24'd239463;
      10'd927: data = 24'd239463;
      10'd928: data = 24'd239463;
      10'd929: data = 24'd239463;
      10'd930: data = 24'd239463;
      10'd931: data = 24'd239463;
      10'd932: data = 24'd239463;
      10'd933: data = 24'd239463;
      10'd934: data = 24'd239463;
      10'd935: data = 24'd239463;
      10'd936: data = 24'd239463;
      10'd937: data = 24'd239463;
      10'd938: data = 24'd239463;
      10'd939: data = 24'd239463;
      10'd940: data = 24'd239463;
      10'd941: data = 24'd239463;
      10'd942: data = 24'd239463;
      10'd943: data = 24'd239463;
      10'd944: data = 24'd239463;
      10'd945: data = 24'd239463;
      10'd946: data = 24'd239463;
      10'd947: data = 24'd239463;
      10'd948: data = 24'd239463;
      10'd949: data = 24'd239463;
      10'd950: data = 24'd239463;
      10'd951: data = 24'd239463;
      10'd952: data = 24'd0;
      10'd953: data = 24'd0;
      10'd954: data = 24'd0;
      10'd955: data = 24'd0;
      10'd956: data = 24'd0;
      10'd957: data = 24'd0;
      10'd958: data = 24'd0;
      10'd959: data = 24'd0;
      10'd960: data = 24'd0;
      10'd961: data = 24'd0;
      10'd962: data = 24'd0;
      10'd963: data = 24'd0;
      10'd964: data = 24'd0;
      10'd965: data = 24'd0;
      10'd966: data = 24'd0;
      10'd967: data = 24'd0;
      10'd968: data = 24'd0;
      10'd969: data = 24'd0;
      10'd970: data = 24'd0;
      10'd971: data = 24'd0;
      10'd972: data = 24'd0;
      10'd973: data = 24'd0;
      10'd974: data = 24'd0;
      10'd975: data = 24'd0;
      10'd976: data = 24'd0;
      10'd977: data = 24'd0;
      10'd978: data = 24'd0;
      10'd979: data = 24'd0;
      10'd980: data = 24'd0;
      10'd981: data = 24'd0;
      10'd982: data = 24'd0;
      10'd983: data = 24'd0;
      10'd984: data = 24'd0;
      10'd985: data = 24'd0;
      10'd986: data = 24'd0;
      10'd987: data = 24'd0;
      10'd988: data = 24'd0;
      10'd989: data = 24'd0;
      10'd990: data = 24'd0;
      10'd991: data = 24'd0;
      10'd992: data = 24'd0;
      10'd993: data = 24'd0;
      10'd994: data = 24'd0;
      10'd995: data = 24'd0;
      10'd996: data = 24'd0;
      10'd997: data = 24'd0;
      10'd998: data = 24'd0;
      10'd999: data = 24'd0;
      10'd1000: data = 24'd0;
      10'd1001: data = 24'd0;
      10'd1002: data = 24'd0;
      10'd1003: data = 24'd0;
      10'd1004: data = 24'd0;
      10'd1005: data = 24'd0;
      10'd1006: data = 24'd0;
      10'd1007: data = 24'd0;
      10'd1008: data = 24'd0;
      10'd1009: data = 24'd0;
      10'd1010: data = 24'd0;
      10'd1011: data = 24'd0;
      10'd1012: data = 24'd0;
      10'd1013: data = 24'd0;
      10'd1014: data = 24'd0;
      10'd1015: data = 24'd0;
      10'd1016: data = 24'd0;
      10'd1017: data = 24'd0;
      10'd1018: data = 24'd0;
      10'd1019: data = 24'd0;
      10'd1020: data = 24'd0;
      10'd1021: data = 24'd0;
      10'd1022: data = 24'd0;
      10'd1023: data = 24'd0;
    endcase
  end
endmodule
